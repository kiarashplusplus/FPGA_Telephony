library verilog;
use verilog.vl_types.all;
entity sys_tb is
end sys_tb;
