library verilog;
use verilog.vl_types.all;
entity combinedTransport_tb is
end combinedTransport_tb;
