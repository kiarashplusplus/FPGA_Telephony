library verilog;
use verilog.vl_types.all;
entity ui_voicemail_test is
end ui_voicemail_test;
